module fmc_top(
    input wire          clk_i,
    input wire          rst_i,

    input wire [24:0]   fmc_a_i,
    input wire          fmc_ne_i,
    input wire          fmc_noe_i,
    input wire          fmc_nwe_i,
    inout      [15:0]   fmc_d_io,
    
    input      [15:0]   fpga_arm_data_i [0:99],
    output     [15:0]   arm_fpga_data_o [0:99]
);
    wire                cs_n;
    wire                rd_n;
    wire                wr_n;
    wire [24:0]         addr;
    wire [15:0]         data;
    wire                noe_tri_en;
    wire [15:0]         fmc_d_o;
    wire [15:0]         fmc_d_i
    assign fmc_noe_i = noe_tri_en?fmc_d_o:16'bzzzz;
    assign fmc_d_i   = fmc_d_io;
    
    fmc_ne_sync fmc_ne_sync_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .fmc_ne_i(fmc_ne_i),
        .cs_o(cs_n)
    );

    fmc_noe_sync fmc_noe_sync_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .fmc_noe_i(fmc_noe_i),
        .rd_o(rd_n)
    );

    fmc_nwe_sync fmc_nwe_sync_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .fmc_nwe_i(fmc_nwe_i),
        .wr_o(wr_n)
    );

    fmc_a_sync fmc_a_sync_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .fmc_a_i(fmc_a_i),
        .addr_o(addr)
    );

    fmc_d_sync fmc_d_sync_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .fmc_d_i(fmc_d_i),
        .data_o(data)
    );
    
    fmc_wr_ram_map fmc_wr_ram_map_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .cs_i(cs_n),
        .rd_i(rd_n),
        .wr_i(wr_n),
        .addr_i(addr),
        .data_i(data),
        .arm_fpga_data_o[0](),
        .arm_fpga_data_o[1](),
        .arm_fpga_data_o[2](),
        .arm_fpga_data_o[3](),
        .arm_fpga_data_o[4](),
        .arm_fpga_data_o[5](),
        .arm_fpga_data_o[6](),
        .arm_fpga_data_o[7](),
        .arm_fpga_data_o[8](),
        .arm_fpga_data_o[9](),
        .arm_fpga_data_o[10](),
        .arm_fpga_data_o[11](),
        .arm_fpga_data_o[12](),
        .arm_fpga_data_o[13](),
        .arm_fpga_data_o[14](),
        .arm_fpga_data_o[15](),
        .arm_fpga_data_o[16](),
        .arm_fpga_data_o[17](),
        .arm_fpga_data_o[18](),
        .arm_fpga_data_o[19](),
        .arm_fpga_data_o[20](),
        .arm_fpga_data_o[21](),
        .arm_fpga_data_o[22](),
        .arm_fpga_data_o[23](),
        .arm_fpga_data_o[24](),
        .arm_fpga_data_o[25](),
        .arm_fpga_data_o[26](),
        .arm_fpga_data_o[27](),
        .arm_fpga_data_o[28](),
        .arm_fpga_data_o[29](),
        .arm_fpga_data_o[30](),
        .arm_fpga_data_o[31](),
        .arm_fpga_data_o[32](),
        .arm_fpga_data_o[33](),
        .arm_fpga_data_o[34](),
        .arm_fpga_data_o[35](),
        .arm_fpga_data_o[36](),
        .arm_fpga_data_o[37](),
        .arm_fpga_data_o[38](),
        .arm_fpga_data_o[39](),
        .arm_fpga_data_o[40](),
        .arm_fpga_data_o[41](),
        .arm_fpga_data_o[42](),
        .arm_fpga_data_o[43](),
        .arm_fpga_data_o[44](),
        .arm_fpga_data_o[45](),
        .arm_fpga_data_o[46](),
        .arm_fpga_data_o[47](),
        .arm_fpga_data_o[48](),
        .arm_fpga_data_o[49](),
        .arm_fpga_data_o[50](),
        .arm_fpga_data_o[51](),
        .arm_fpga_data_o[52](),
        .arm_fpga_data_o[53](),
        .arm_fpga_data_o[54](),
        .arm_fpga_data_o[55](),
        .arm_fpga_data_o[56](),
        .arm_fpga_data_o[57](),
        .arm_fpga_data_o[58](),
        .arm_fpga_data_o[59](),
        .arm_fpga_data_o[60](),
        .arm_fpga_data_o[61](),
        .arm_fpga_data_o[62](),
        .arm_fpga_data_o[63](),
        .arm_fpga_data_o[64](),
        .arm_fpga_data_o[65](),
        .arm_fpga_data_o[66](),
        .arm_fpga_data_o[67](),
        .arm_fpga_data_o[68](),
        .arm_fpga_data_o[69](),
        .arm_fpga_data_o[70](),
        .arm_fpga_data_o[71](),
        .arm_fpga_data_o[72](),
        .arm_fpga_data_o[73](),
        .arm_fpga_data_o[74](),
        .arm_fpga_data_o[75](),
        .arm_fpga_data_o[76](),
        .arm_fpga_data_o[77](),
        .arm_fpga_data_o[78](),
        .arm_fpga_data_o[79](),
        .arm_fpga_data_o[80](),
        .arm_fpga_data_o[81](),
        .arm_fpga_data_o[82](),
        .arm_fpga_data_o[83](),
        .arm_fpga_data_o[84](),
        .arm_fpga_data_o[85](),
        .arm_fpga_data_o[86](),
        .arm_fpga_data_o[87](),
        .arm_fpga_data_o[88](),
        .arm_fpga_data_o[89](),
        .arm_fpga_data_o[90](),
        .arm_fpga_data_o[91](),
        .arm_fpga_data_o[92](),
        .arm_fpga_data_o[93](),
        .arm_fpga_data_o[94](),
        .arm_fpga_data_o[95](),
        .arm_fpga_data_o[96](),
        .arm_fpga_data_o[97](),
        .arm_fpga_data_o[98](),
        .arm_fpga_data_o[99]()
    );

    fmc_rd_ram_map fmc_rd_ram_map_init(
        .clk_i(clk_i),
        .rst_i(rst_i),
        .cs_i(cs_n),
        .rd_i(rd_n),
        .wr_i(wr_n),
        .addr_i(addr),
        .thr_state_en(noe_tri_en),
        .data_o(fmc_d_o),
        .fpga_arm_data_i[0](),
        .fpga_arm_data_i[1](),
        .fpga_arm_data_i[2](),
        .fpga_arm_data_i[3](),
        .fpga_arm_data_i[4](),
        .fpga_arm_data_i[5](),
        .fpga_arm_data_i[6](),
        .fpga_arm_data_i[7](),
        .fpga_arm_data_i[8](),
        .fpga_arm_data_i[9](),
        .fpga_arm_data_i[10](),
        .fpga_arm_data_i[11](),
        .fpga_arm_data_i[12](),
        .fpga_arm_data_i[13](),
        .fpga_arm_data_i[14](),
        .fpga_arm_data_i[15](),
        .fpga_arm_data_i[16](),
        .fpga_arm_data_i[17](),
        .fpga_arm_data_i[18](),
        .fpga_arm_data_i[19](),
        .fpga_arm_data_i[20](),
        .fpga_arm_data_i[21](),
        .fpga_arm_data_i[22](),
        .fpga_arm_data_i[23](),
        .fpga_arm_data_i[24](),
        .fpga_arm_data_i[25](),
        .fpga_arm_data_i[26](),
        .fpga_arm_data_i[27](),
        .fpga_arm_data_i[28](),
        .fpga_arm_data_i[29](),
        .fpga_arm_data_i[30](),
        .fpga_arm_data_i[31](),
        .fpga_arm_data_i[32](),
        .fpga_arm_data_i[33](),
        .fpga_arm_data_i[34](),
        .fpga_arm_data_i[35](),
        .fpga_arm_data_i[36](),
        .fpga_arm_data_i[37](),
        .fpga_arm_data_i[38](),
        .fpga_arm_data_i[39](),
        .fpga_arm_data_i[40](),
        .fpga_arm_data_i[41](),
        .fpga_arm_data_i[42](),
        .fpga_arm_data_i[43](),
        .fpga_arm_data_i[44](),
        .fpga_arm_data_i[45](),
        .fpga_arm_data_i[46](),
        .fpga_arm_data_i[47](),
        .fpga_arm_data_i[48](),
        .fpga_arm_data_i[49](),
        .fpga_arm_data_i[50](),
        .fpga_arm_data_i[51](),
        .fpga_arm_data_i[52](),
        .fpga_arm_data_i[53](),
        .fpga_arm_data_i[54](),
        .fpga_arm_data_i[55](),
        .fpga_arm_data_i[56](),
        .fpga_arm_data_i[57](),
        .fpga_arm_data_i[58](),
        .fpga_arm_data_i[59](),
        .fpga_arm_data_i[60](),
        .fpga_arm_data_i[61](),
        .fpga_arm_data_i[62](),
        .fpga_arm_data_i[63](),
        .fpga_arm_data_i[64](),
        .fpga_arm_data_i[65](),
        .fpga_arm_data_i[66](),
        .fpga_arm_data_i[67](),
        .fpga_arm_data_i[68](),
        .fpga_arm_data_i[69](),
        .fpga_arm_data_i[70](),
        .fpga_arm_data_i[71](),
        .fpga_arm_data_i[72](),
        .fpga_arm_data_i[73](),
        .fpga_arm_data_i[74](),
        .fpga_arm_data_i[75](),
        .fpga_arm_data_i[76](),
        .fpga_arm_data_i[77](),
        .fpga_arm_data_i[78](),
        .fpga_arm_data_i[79](),
        .fpga_arm_data_i[80](),
        .fpga_arm_data_i[81](),
        .fpga_arm_data_i[82](),
        .fpga_arm_data_i[83](),
        .fpga_arm_data_i[84](),
        .fpga_arm_data_i[85](),
        .fpga_arm_data_i[86](),
        .fpga_arm_data_i[87](),
        .fpga_arm_data_i[88](),
        .fpga_arm_data_i[89](),
        .fpga_arm_data_i[90](),
        .fpga_arm_data_i[91](),
        .fpga_arm_data_i[92](),
        .fpga_arm_data_i[93](),
        .fpga_arm_data_i[94](),
        .fpga_arm_data_i[95](),
        .fpga_arm_data_i[96](),
        .fpga_arm_data_i[97](),
        .fpga_arm_data_i[98](),
        .fpga_arm_data_i[99]()
    );


endmodule